module gw_gao(
    \read_data[15] ,
    \read_data[14] ,
    \read_data[13] ,
    \read_data[12] ,
    \read_data[11] ,
    \read_data[10] ,
    \read_data[9] ,
    \read_data[8] ,
    \read_data[7] ,
    \read_data[6] ,
    \read_data[5] ,
    \read_data[4] ,
    \read_data[3] ,
    \read_data[2] ,
    \read_data[1] ,
    \read_data[0] ,
    \fifo_ram_module/rd_data[255] ,
    \fifo_ram_module/rd_data[254] ,
    \fifo_ram_module/rd_data[253] ,
    \fifo_ram_module/rd_data[252] ,
    \fifo_ram_module/rd_data[251] ,
    \fifo_ram_module/rd_data[250] ,
    \fifo_ram_module/rd_data[249] ,
    \fifo_ram_module/rd_data[248] ,
    \fifo_ram_module/rd_data[247] ,
    \fifo_ram_module/rd_data[246] ,
    \fifo_ram_module/rd_data[245] ,
    \fifo_ram_module/rd_data[244] ,
    \fifo_ram_module/rd_data[243] ,
    \fifo_ram_module/rd_data[242] ,
    \fifo_ram_module/rd_data[241] ,
    \fifo_ram_module/rd_data[240] ,
    \fifo_ram_module/rd_data[239] ,
    \fifo_ram_module/rd_data[238] ,
    \fifo_ram_module/rd_data[237] ,
    \fifo_ram_module/rd_data[236] ,
    \fifo_ram_module/rd_data[235] ,
    \fifo_ram_module/rd_data[234] ,
    \fifo_ram_module/rd_data[233] ,
    \fifo_ram_module/rd_data[232] ,
    \fifo_ram_module/rd_data[231] ,
    \fifo_ram_module/rd_data[230] ,
    \fifo_ram_module/rd_data[229] ,
    \fifo_ram_module/rd_data[228] ,
    \fifo_ram_module/rd_data[227] ,
    \fifo_ram_module/rd_data[226] ,
    \fifo_ram_module/rd_data[225] ,
    \fifo_ram_module/rd_data[224] ,
    \fifo_ram_module/rd_data[223] ,
    \fifo_ram_module/rd_data[222] ,
    \fifo_ram_module/rd_data[221] ,
    \fifo_ram_module/rd_data[220] ,
    \fifo_ram_module/rd_data[219] ,
    \fifo_ram_module/rd_data[218] ,
    \fifo_ram_module/rd_data[217] ,
    \fifo_ram_module/rd_data[216] ,
    \fifo_ram_module/rd_data[215] ,
    \fifo_ram_module/rd_data[214] ,
    \fifo_ram_module/rd_data[213] ,
    \fifo_ram_module/rd_data[212] ,
    \fifo_ram_module/rd_data[211] ,
    \fifo_ram_module/rd_data[210] ,
    \fifo_ram_module/rd_data[209] ,
    \fifo_ram_module/rd_data[208] ,
    \fifo_ram_module/rd_data[207] ,
    \fifo_ram_module/rd_data[206] ,
    \fifo_ram_module/rd_data[205] ,
    \fifo_ram_module/rd_data[204] ,
    \fifo_ram_module/rd_data[203] ,
    \fifo_ram_module/rd_data[202] ,
    \fifo_ram_module/rd_data[201] ,
    \fifo_ram_module/rd_data[200] ,
    \fifo_ram_module/rd_data[199] ,
    \fifo_ram_module/rd_data[198] ,
    \fifo_ram_module/rd_data[197] ,
    \fifo_ram_module/rd_data[196] ,
    \fifo_ram_module/rd_data[195] ,
    \fifo_ram_module/rd_data[194] ,
    \fifo_ram_module/rd_data[193] ,
    \fifo_ram_module/rd_data[192] ,
    \fifo_ram_module/rd_data[191] ,
    \fifo_ram_module/rd_data[190] ,
    \fifo_ram_module/rd_data[189] ,
    \fifo_ram_module/rd_data[188] ,
    \fifo_ram_module/rd_data[187] ,
    \fifo_ram_module/rd_data[186] ,
    \fifo_ram_module/rd_data[185] ,
    \fifo_ram_module/rd_data[184] ,
    \fifo_ram_module/rd_data[183] ,
    \fifo_ram_module/rd_data[182] ,
    \fifo_ram_module/rd_data[181] ,
    \fifo_ram_module/rd_data[180] ,
    \fifo_ram_module/rd_data[179] ,
    \fifo_ram_module/rd_data[178] ,
    \fifo_ram_module/rd_data[177] ,
    \fifo_ram_module/rd_data[176] ,
    \fifo_ram_module/rd_data[175] ,
    \fifo_ram_module/rd_data[174] ,
    \fifo_ram_module/rd_data[173] ,
    \fifo_ram_module/rd_data[172] ,
    \fifo_ram_module/rd_data[171] ,
    \fifo_ram_module/rd_data[170] ,
    \fifo_ram_module/rd_data[169] ,
    \fifo_ram_module/rd_data[168] ,
    \fifo_ram_module/rd_data[167] ,
    \fifo_ram_module/rd_data[166] ,
    \fifo_ram_module/rd_data[165] ,
    \fifo_ram_module/rd_data[164] ,
    \fifo_ram_module/rd_data[163] ,
    \fifo_ram_module/rd_data[162] ,
    \fifo_ram_module/rd_data[161] ,
    \fifo_ram_module/rd_data[160] ,
    \fifo_ram_module/rd_data[159] ,
    \fifo_ram_module/rd_data[158] ,
    \fifo_ram_module/rd_data[157] ,
    \fifo_ram_module/rd_data[156] ,
    \fifo_ram_module/rd_data[155] ,
    \fifo_ram_module/rd_data[154] ,
    \fifo_ram_module/rd_data[153] ,
    \fifo_ram_module/rd_data[152] ,
    \fifo_ram_module/rd_data[151] ,
    \fifo_ram_module/rd_data[150] ,
    \fifo_ram_module/rd_data[149] ,
    \fifo_ram_module/rd_data[148] ,
    \fifo_ram_module/rd_data[147] ,
    \fifo_ram_module/rd_data[146] ,
    \fifo_ram_module/rd_data[145] ,
    \fifo_ram_module/rd_data[144] ,
    \fifo_ram_module/rd_data[143] ,
    \fifo_ram_module/rd_data[142] ,
    \fifo_ram_module/rd_data[141] ,
    \fifo_ram_module/rd_data[140] ,
    \fifo_ram_module/rd_data[139] ,
    \fifo_ram_module/rd_data[138] ,
    \fifo_ram_module/rd_data[137] ,
    \fifo_ram_module/rd_data[136] ,
    \fifo_ram_module/rd_data[135] ,
    \fifo_ram_module/rd_data[134] ,
    \fifo_ram_module/rd_data[133] ,
    \fifo_ram_module/rd_data[132] ,
    \fifo_ram_module/rd_data[131] ,
    \fifo_ram_module/rd_data[130] ,
    \fifo_ram_module/rd_data[129] ,
    \fifo_ram_module/rd_data[128] ,
    \fifo_ram_module/rd_data[127] ,
    \fifo_ram_module/rd_data[126] ,
    \fifo_ram_module/rd_data[125] ,
    \fifo_ram_module/rd_data[124] ,
    \fifo_ram_module/rd_data[123] ,
    \fifo_ram_module/rd_data[122] ,
    \fifo_ram_module/rd_data[121] ,
    \fifo_ram_module/rd_data[120] ,
    \fifo_ram_module/rd_data[119] ,
    \fifo_ram_module/rd_data[118] ,
    \fifo_ram_module/rd_data[117] ,
    \fifo_ram_module/rd_data[116] ,
    \fifo_ram_module/rd_data[115] ,
    \fifo_ram_module/rd_data[114] ,
    \fifo_ram_module/rd_data[113] ,
    \fifo_ram_module/rd_data[112] ,
    \fifo_ram_module/rd_data[111] ,
    \fifo_ram_module/rd_data[110] ,
    \fifo_ram_module/rd_data[109] ,
    \fifo_ram_module/rd_data[108] ,
    \fifo_ram_module/rd_data[107] ,
    \fifo_ram_module/rd_data[106] ,
    \fifo_ram_module/rd_data[105] ,
    \fifo_ram_module/rd_data[104] ,
    \fifo_ram_module/rd_data[103] ,
    \fifo_ram_module/rd_data[102] ,
    \fifo_ram_module/rd_data[101] ,
    \fifo_ram_module/rd_data[100] ,
    \fifo_ram_module/rd_data[99] ,
    \fifo_ram_module/rd_data[98] ,
    \fifo_ram_module/rd_data[97] ,
    \fifo_ram_module/rd_data[96] ,
    \fifo_ram_module/rd_data[95] ,
    \fifo_ram_module/rd_data[94] ,
    \fifo_ram_module/rd_data[93] ,
    \fifo_ram_module/rd_data[92] ,
    \fifo_ram_module/rd_data[91] ,
    \fifo_ram_module/rd_data[90] ,
    \fifo_ram_module/rd_data[89] ,
    \fifo_ram_module/rd_data[88] ,
    \fifo_ram_module/rd_data[87] ,
    \fifo_ram_module/rd_data[86] ,
    \fifo_ram_module/rd_data[85] ,
    \fifo_ram_module/rd_data[84] ,
    \fifo_ram_module/rd_data[83] ,
    \fifo_ram_module/rd_data[82] ,
    \fifo_ram_module/rd_data[81] ,
    \fifo_ram_module/rd_data[80] ,
    \fifo_ram_module/rd_data[79] ,
    \fifo_ram_module/rd_data[78] ,
    \fifo_ram_module/rd_data[77] ,
    \fifo_ram_module/rd_data[76] ,
    \fifo_ram_module/rd_data[75] ,
    \fifo_ram_module/rd_data[74] ,
    \fifo_ram_module/rd_data[73] ,
    \fifo_ram_module/rd_data[72] ,
    \fifo_ram_module/rd_data[71] ,
    \fifo_ram_module/rd_data[70] ,
    \fifo_ram_module/rd_data[69] ,
    \fifo_ram_module/rd_data[68] ,
    \fifo_ram_module/rd_data[67] ,
    \fifo_ram_module/rd_data[66] ,
    \fifo_ram_module/rd_data[65] ,
    \fifo_ram_module/rd_data[64] ,
    \fifo_ram_module/rd_data[63] ,
    \fifo_ram_module/rd_data[62] ,
    \fifo_ram_module/rd_data[61] ,
    \fifo_ram_module/rd_data[60] ,
    \fifo_ram_module/rd_data[59] ,
    \fifo_ram_module/rd_data[58] ,
    \fifo_ram_module/rd_data[57] ,
    \fifo_ram_module/rd_data[56] ,
    \fifo_ram_module/rd_data[55] ,
    \fifo_ram_module/rd_data[54] ,
    \fifo_ram_module/rd_data[53] ,
    \fifo_ram_module/rd_data[52] ,
    \fifo_ram_module/rd_data[51] ,
    \fifo_ram_module/rd_data[50] ,
    \fifo_ram_module/rd_data[49] ,
    \fifo_ram_module/rd_data[48] ,
    \fifo_ram_module/rd_data[47] ,
    \fifo_ram_module/rd_data[46] ,
    \fifo_ram_module/rd_data[45] ,
    \fifo_ram_module/rd_data[44] ,
    \fifo_ram_module/rd_data[43] ,
    \fifo_ram_module/rd_data[42] ,
    \fifo_ram_module/rd_data[41] ,
    \fifo_ram_module/rd_data[40] ,
    \fifo_ram_module/rd_data[39] ,
    \fifo_ram_module/rd_data[38] ,
    \fifo_ram_module/rd_data[37] ,
    \fifo_ram_module/rd_data[36] ,
    \fifo_ram_module/rd_data[35] ,
    \fifo_ram_module/rd_data[34] ,
    \fifo_ram_module/rd_data[33] ,
    \fifo_ram_module/rd_data[32] ,
    \fifo_ram_module/rd_data[31] ,
    \fifo_ram_module/rd_data[30] ,
    \fifo_ram_module/rd_data[29] ,
    \fifo_ram_module/rd_data[28] ,
    \fifo_ram_module/rd_data[27] ,
    \fifo_ram_module/rd_data[26] ,
    \fifo_ram_module/rd_data[25] ,
    \fifo_ram_module/rd_data[24] ,
    \fifo_ram_module/rd_data[23] ,
    \fifo_ram_module/rd_data[22] ,
    \fifo_ram_module/rd_data[21] ,
    \fifo_ram_module/rd_data[20] ,
    \fifo_ram_module/rd_data[19] ,
    \fifo_ram_module/rd_data[18] ,
    \fifo_ram_module/rd_data[17] ,
    \fifo_ram_module/rd_data[16] ,
    \fifo_ram_module/rd_data[15] ,
    \fifo_ram_module/rd_data[14] ,
    \fifo_ram_module/rd_data[13] ,
    \fifo_ram_module/rd_data[12] ,
    \fifo_ram_module/rd_data[11] ,
    \fifo_ram_module/rd_data[10] ,
    \fifo_ram_module/rd_data[9] ,
    \fifo_ram_module/rd_data[8] ,
    \fifo_ram_module/rd_data[7] ,
    \fifo_ram_module/rd_data[6] ,
    \fifo_ram_module/rd_data[5] ,
    \fifo_ram_module/rd_data[4] ,
    \fifo_ram_module/rd_data[3] ,
    \fifo_ram_module/rd_data[2] ,
    \fifo_ram_module/rd_data[1] ,
    \fifo_ram_module/rd_data[0] ,
    \fifo_ram_module/cmd[2] ,
    \fifo_ram_module/cmd[1] ,
    \fifo_ram_module/cmd[0] ,
    \fifo_ram_module/app_addr[28] ,
    \fifo_ram_module/app_addr[27] ,
    \fifo_ram_module/app_addr[26] ,
    \fifo_ram_module/app_addr[25] ,
    \fifo_ram_module/app_addr[24] ,
    \fifo_ram_module/app_addr[23] ,
    \fifo_ram_module/app_addr[22] ,
    \fifo_ram_module/app_addr[21] ,
    \fifo_ram_module/app_addr[20] ,
    \fifo_ram_module/app_addr[19] ,
    \fifo_ram_module/app_addr[18] ,
    \fifo_ram_module/app_addr[17] ,
    \fifo_ram_module/app_addr[16] ,
    \fifo_ram_module/app_addr[15] ,
    \fifo_ram_module/app_addr[14] ,
    \fifo_ram_module/app_addr[13] ,
    \fifo_ram_module/app_addr[12] ,
    \fifo_ram_module/app_addr[11] ,
    \fifo_ram_module/app_addr[10] ,
    \fifo_ram_module/app_addr[9] ,
    \fifo_ram_module/app_addr[8] ,
    \fifo_ram_module/app_addr[7] ,
    \fifo_ram_module/app_addr[6] ,
    \fifo_ram_module/app_addr[5] ,
    \fifo_ram_module/app_addr[4] ,
    \fifo_ram_module/app_addr[3] ,
    \fifo_ram_module/app_addr[2] ,
    \fifo_ram_module/app_addr[1] ,
    \fifo_ram_module/app_addr[0] ,
    \fifo_ram_module/state[3] ,
    \fifo_ram_module/state[2] ,
    \fifo_ram_module/state[1] ,
    \fifo_ram_module/state[0] ,
    \fifo_ram_module/count[31] ,
    \fifo_ram_module/count[30] ,
    \fifo_ram_module/count[29] ,
    \fifo_ram_module/count[28] ,
    \fifo_ram_module/count[27] ,
    \fifo_ram_module/count[26] ,
    \fifo_ram_module/count[25] ,
    \fifo_ram_module/count[24] ,
    \fifo_ram_module/count[23] ,
    \fifo_ram_module/count[22] ,
    \fifo_ram_module/count[21] ,
    \fifo_ram_module/count[20] ,
    \fifo_ram_module/count[19] ,
    \fifo_ram_module/count[18] ,
    \fifo_ram_module/count[17] ,
    \fifo_ram_module/count[16] ,
    \fifo_ram_module/count[15] ,
    \fifo_ram_module/count[14] ,
    \fifo_ram_module/count[13] ,
    \fifo_ram_module/count[12] ,
    \fifo_ram_module/count[11] ,
    \fifo_ram_module/count[10] ,
    \fifo_ram_module/count[9] ,
    \fifo_ram_module/count[8] ,
    \fifo_ram_module/count[7] ,
    \fifo_ram_module/count[6] ,
    \fifo_ram_module/count[5] ,
    \fifo_ram_module/count[4] ,
    \fifo_ram_module/count[3] ,
    \fifo_ram_module/count[2] ,
    \fifo_ram_module/count[1] ,
    \fifo_ram_module/count[0] ,
    \fifo_ram_module/cmd_ready ,
    \fifo_ram_module/cmd_en ,
    \fifo_ram_module/wr_ready ,
    \fifo_ram_module/wr_en ,
    \fifo_ram_module/rd_data_valid ,
    \fifo_ram_module/fifo_read_full ,
    \fifo_ram_module/fifo_write_empty ,
    \fifo_ram_module/fifo_read_almost_empty ,
    \fifo_ram_module/fifo_write_rd_en ,
    \fifo_ram_module/fifo_read_wr_en ,
    \fifo_ram_module/fifo_write_full ,
    \fifo_ram_module/fifo_read_empty ,
    read_en,
    \state[3] ,
    \state[2] ,
    \state[1] ,
    \state[0] ,
    sd_file_found,
    clk,
    tms_pad_i,
    tck_pad_i,
    tdi_pad_i,
    tdo_pad_o
);

input \read_data[15] ;
input \read_data[14] ;
input \read_data[13] ;
input \read_data[12] ;
input \read_data[11] ;
input \read_data[10] ;
input \read_data[9] ;
input \read_data[8] ;
input \read_data[7] ;
input \read_data[6] ;
input \read_data[5] ;
input \read_data[4] ;
input \read_data[3] ;
input \read_data[2] ;
input \read_data[1] ;
input \read_data[0] ;
input \fifo_ram_module/rd_data[255] ;
input \fifo_ram_module/rd_data[254] ;
input \fifo_ram_module/rd_data[253] ;
input \fifo_ram_module/rd_data[252] ;
input \fifo_ram_module/rd_data[251] ;
input \fifo_ram_module/rd_data[250] ;
input \fifo_ram_module/rd_data[249] ;
input \fifo_ram_module/rd_data[248] ;
input \fifo_ram_module/rd_data[247] ;
input \fifo_ram_module/rd_data[246] ;
input \fifo_ram_module/rd_data[245] ;
input \fifo_ram_module/rd_data[244] ;
input \fifo_ram_module/rd_data[243] ;
input \fifo_ram_module/rd_data[242] ;
input \fifo_ram_module/rd_data[241] ;
input \fifo_ram_module/rd_data[240] ;
input \fifo_ram_module/rd_data[239] ;
input \fifo_ram_module/rd_data[238] ;
input \fifo_ram_module/rd_data[237] ;
input \fifo_ram_module/rd_data[236] ;
input \fifo_ram_module/rd_data[235] ;
input \fifo_ram_module/rd_data[234] ;
input \fifo_ram_module/rd_data[233] ;
input \fifo_ram_module/rd_data[232] ;
input \fifo_ram_module/rd_data[231] ;
input \fifo_ram_module/rd_data[230] ;
input \fifo_ram_module/rd_data[229] ;
input \fifo_ram_module/rd_data[228] ;
input \fifo_ram_module/rd_data[227] ;
input \fifo_ram_module/rd_data[226] ;
input \fifo_ram_module/rd_data[225] ;
input \fifo_ram_module/rd_data[224] ;
input \fifo_ram_module/rd_data[223] ;
input \fifo_ram_module/rd_data[222] ;
input \fifo_ram_module/rd_data[221] ;
input \fifo_ram_module/rd_data[220] ;
input \fifo_ram_module/rd_data[219] ;
input \fifo_ram_module/rd_data[218] ;
input \fifo_ram_module/rd_data[217] ;
input \fifo_ram_module/rd_data[216] ;
input \fifo_ram_module/rd_data[215] ;
input \fifo_ram_module/rd_data[214] ;
input \fifo_ram_module/rd_data[213] ;
input \fifo_ram_module/rd_data[212] ;
input \fifo_ram_module/rd_data[211] ;
input \fifo_ram_module/rd_data[210] ;
input \fifo_ram_module/rd_data[209] ;
input \fifo_ram_module/rd_data[208] ;
input \fifo_ram_module/rd_data[207] ;
input \fifo_ram_module/rd_data[206] ;
input \fifo_ram_module/rd_data[205] ;
input \fifo_ram_module/rd_data[204] ;
input \fifo_ram_module/rd_data[203] ;
input \fifo_ram_module/rd_data[202] ;
input \fifo_ram_module/rd_data[201] ;
input \fifo_ram_module/rd_data[200] ;
input \fifo_ram_module/rd_data[199] ;
input \fifo_ram_module/rd_data[198] ;
input \fifo_ram_module/rd_data[197] ;
input \fifo_ram_module/rd_data[196] ;
input \fifo_ram_module/rd_data[195] ;
input \fifo_ram_module/rd_data[194] ;
input \fifo_ram_module/rd_data[193] ;
input \fifo_ram_module/rd_data[192] ;
input \fifo_ram_module/rd_data[191] ;
input \fifo_ram_module/rd_data[190] ;
input \fifo_ram_module/rd_data[189] ;
input \fifo_ram_module/rd_data[188] ;
input \fifo_ram_module/rd_data[187] ;
input \fifo_ram_module/rd_data[186] ;
input \fifo_ram_module/rd_data[185] ;
input \fifo_ram_module/rd_data[184] ;
input \fifo_ram_module/rd_data[183] ;
input \fifo_ram_module/rd_data[182] ;
input \fifo_ram_module/rd_data[181] ;
input \fifo_ram_module/rd_data[180] ;
input \fifo_ram_module/rd_data[179] ;
input \fifo_ram_module/rd_data[178] ;
input \fifo_ram_module/rd_data[177] ;
input \fifo_ram_module/rd_data[176] ;
input \fifo_ram_module/rd_data[175] ;
input \fifo_ram_module/rd_data[174] ;
input \fifo_ram_module/rd_data[173] ;
input \fifo_ram_module/rd_data[172] ;
input \fifo_ram_module/rd_data[171] ;
input \fifo_ram_module/rd_data[170] ;
input \fifo_ram_module/rd_data[169] ;
input \fifo_ram_module/rd_data[168] ;
input \fifo_ram_module/rd_data[167] ;
input \fifo_ram_module/rd_data[166] ;
input \fifo_ram_module/rd_data[165] ;
input \fifo_ram_module/rd_data[164] ;
input \fifo_ram_module/rd_data[163] ;
input \fifo_ram_module/rd_data[162] ;
input \fifo_ram_module/rd_data[161] ;
input \fifo_ram_module/rd_data[160] ;
input \fifo_ram_module/rd_data[159] ;
input \fifo_ram_module/rd_data[158] ;
input \fifo_ram_module/rd_data[157] ;
input \fifo_ram_module/rd_data[156] ;
input \fifo_ram_module/rd_data[155] ;
input \fifo_ram_module/rd_data[154] ;
input \fifo_ram_module/rd_data[153] ;
input \fifo_ram_module/rd_data[152] ;
input \fifo_ram_module/rd_data[151] ;
input \fifo_ram_module/rd_data[150] ;
input \fifo_ram_module/rd_data[149] ;
input \fifo_ram_module/rd_data[148] ;
input \fifo_ram_module/rd_data[147] ;
input \fifo_ram_module/rd_data[146] ;
input \fifo_ram_module/rd_data[145] ;
input \fifo_ram_module/rd_data[144] ;
input \fifo_ram_module/rd_data[143] ;
input \fifo_ram_module/rd_data[142] ;
input \fifo_ram_module/rd_data[141] ;
input \fifo_ram_module/rd_data[140] ;
input \fifo_ram_module/rd_data[139] ;
input \fifo_ram_module/rd_data[138] ;
input \fifo_ram_module/rd_data[137] ;
input \fifo_ram_module/rd_data[136] ;
input \fifo_ram_module/rd_data[135] ;
input \fifo_ram_module/rd_data[134] ;
input \fifo_ram_module/rd_data[133] ;
input \fifo_ram_module/rd_data[132] ;
input \fifo_ram_module/rd_data[131] ;
input \fifo_ram_module/rd_data[130] ;
input \fifo_ram_module/rd_data[129] ;
input \fifo_ram_module/rd_data[128] ;
input \fifo_ram_module/rd_data[127] ;
input \fifo_ram_module/rd_data[126] ;
input \fifo_ram_module/rd_data[125] ;
input \fifo_ram_module/rd_data[124] ;
input \fifo_ram_module/rd_data[123] ;
input \fifo_ram_module/rd_data[122] ;
input \fifo_ram_module/rd_data[121] ;
input \fifo_ram_module/rd_data[120] ;
input \fifo_ram_module/rd_data[119] ;
input \fifo_ram_module/rd_data[118] ;
input \fifo_ram_module/rd_data[117] ;
input \fifo_ram_module/rd_data[116] ;
input \fifo_ram_module/rd_data[115] ;
input \fifo_ram_module/rd_data[114] ;
input \fifo_ram_module/rd_data[113] ;
input \fifo_ram_module/rd_data[112] ;
input \fifo_ram_module/rd_data[111] ;
input \fifo_ram_module/rd_data[110] ;
input \fifo_ram_module/rd_data[109] ;
input \fifo_ram_module/rd_data[108] ;
input \fifo_ram_module/rd_data[107] ;
input \fifo_ram_module/rd_data[106] ;
input \fifo_ram_module/rd_data[105] ;
input \fifo_ram_module/rd_data[104] ;
input \fifo_ram_module/rd_data[103] ;
input \fifo_ram_module/rd_data[102] ;
input \fifo_ram_module/rd_data[101] ;
input \fifo_ram_module/rd_data[100] ;
input \fifo_ram_module/rd_data[99] ;
input \fifo_ram_module/rd_data[98] ;
input \fifo_ram_module/rd_data[97] ;
input \fifo_ram_module/rd_data[96] ;
input \fifo_ram_module/rd_data[95] ;
input \fifo_ram_module/rd_data[94] ;
input \fifo_ram_module/rd_data[93] ;
input \fifo_ram_module/rd_data[92] ;
input \fifo_ram_module/rd_data[91] ;
input \fifo_ram_module/rd_data[90] ;
input \fifo_ram_module/rd_data[89] ;
input \fifo_ram_module/rd_data[88] ;
input \fifo_ram_module/rd_data[87] ;
input \fifo_ram_module/rd_data[86] ;
input \fifo_ram_module/rd_data[85] ;
input \fifo_ram_module/rd_data[84] ;
input \fifo_ram_module/rd_data[83] ;
input \fifo_ram_module/rd_data[82] ;
input \fifo_ram_module/rd_data[81] ;
input \fifo_ram_module/rd_data[80] ;
input \fifo_ram_module/rd_data[79] ;
input \fifo_ram_module/rd_data[78] ;
input \fifo_ram_module/rd_data[77] ;
input \fifo_ram_module/rd_data[76] ;
input \fifo_ram_module/rd_data[75] ;
input \fifo_ram_module/rd_data[74] ;
input \fifo_ram_module/rd_data[73] ;
input \fifo_ram_module/rd_data[72] ;
input \fifo_ram_module/rd_data[71] ;
input \fifo_ram_module/rd_data[70] ;
input \fifo_ram_module/rd_data[69] ;
input \fifo_ram_module/rd_data[68] ;
input \fifo_ram_module/rd_data[67] ;
input \fifo_ram_module/rd_data[66] ;
input \fifo_ram_module/rd_data[65] ;
input \fifo_ram_module/rd_data[64] ;
input \fifo_ram_module/rd_data[63] ;
input \fifo_ram_module/rd_data[62] ;
input \fifo_ram_module/rd_data[61] ;
input \fifo_ram_module/rd_data[60] ;
input \fifo_ram_module/rd_data[59] ;
input \fifo_ram_module/rd_data[58] ;
input \fifo_ram_module/rd_data[57] ;
input \fifo_ram_module/rd_data[56] ;
input \fifo_ram_module/rd_data[55] ;
input \fifo_ram_module/rd_data[54] ;
input \fifo_ram_module/rd_data[53] ;
input \fifo_ram_module/rd_data[52] ;
input \fifo_ram_module/rd_data[51] ;
input \fifo_ram_module/rd_data[50] ;
input \fifo_ram_module/rd_data[49] ;
input \fifo_ram_module/rd_data[48] ;
input \fifo_ram_module/rd_data[47] ;
input \fifo_ram_module/rd_data[46] ;
input \fifo_ram_module/rd_data[45] ;
input \fifo_ram_module/rd_data[44] ;
input \fifo_ram_module/rd_data[43] ;
input \fifo_ram_module/rd_data[42] ;
input \fifo_ram_module/rd_data[41] ;
input \fifo_ram_module/rd_data[40] ;
input \fifo_ram_module/rd_data[39] ;
input \fifo_ram_module/rd_data[38] ;
input \fifo_ram_module/rd_data[37] ;
input \fifo_ram_module/rd_data[36] ;
input \fifo_ram_module/rd_data[35] ;
input \fifo_ram_module/rd_data[34] ;
input \fifo_ram_module/rd_data[33] ;
input \fifo_ram_module/rd_data[32] ;
input \fifo_ram_module/rd_data[31] ;
input \fifo_ram_module/rd_data[30] ;
input \fifo_ram_module/rd_data[29] ;
input \fifo_ram_module/rd_data[28] ;
input \fifo_ram_module/rd_data[27] ;
input \fifo_ram_module/rd_data[26] ;
input \fifo_ram_module/rd_data[25] ;
input \fifo_ram_module/rd_data[24] ;
input \fifo_ram_module/rd_data[23] ;
input \fifo_ram_module/rd_data[22] ;
input \fifo_ram_module/rd_data[21] ;
input \fifo_ram_module/rd_data[20] ;
input \fifo_ram_module/rd_data[19] ;
input \fifo_ram_module/rd_data[18] ;
input \fifo_ram_module/rd_data[17] ;
input \fifo_ram_module/rd_data[16] ;
input \fifo_ram_module/rd_data[15] ;
input \fifo_ram_module/rd_data[14] ;
input \fifo_ram_module/rd_data[13] ;
input \fifo_ram_module/rd_data[12] ;
input \fifo_ram_module/rd_data[11] ;
input \fifo_ram_module/rd_data[10] ;
input \fifo_ram_module/rd_data[9] ;
input \fifo_ram_module/rd_data[8] ;
input \fifo_ram_module/rd_data[7] ;
input \fifo_ram_module/rd_data[6] ;
input \fifo_ram_module/rd_data[5] ;
input \fifo_ram_module/rd_data[4] ;
input \fifo_ram_module/rd_data[3] ;
input \fifo_ram_module/rd_data[2] ;
input \fifo_ram_module/rd_data[1] ;
input \fifo_ram_module/rd_data[0] ;
input \fifo_ram_module/cmd[2] ;
input \fifo_ram_module/cmd[1] ;
input \fifo_ram_module/cmd[0] ;
input \fifo_ram_module/app_addr[28] ;
input \fifo_ram_module/app_addr[27] ;
input \fifo_ram_module/app_addr[26] ;
input \fifo_ram_module/app_addr[25] ;
input \fifo_ram_module/app_addr[24] ;
input \fifo_ram_module/app_addr[23] ;
input \fifo_ram_module/app_addr[22] ;
input \fifo_ram_module/app_addr[21] ;
input \fifo_ram_module/app_addr[20] ;
input \fifo_ram_module/app_addr[19] ;
input \fifo_ram_module/app_addr[18] ;
input \fifo_ram_module/app_addr[17] ;
input \fifo_ram_module/app_addr[16] ;
input \fifo_ram_module/app_addr[15] ;
input \fifo_ram_module/app_addr[14] ;
input \fifo_ram_module/app_addr[13] ;
input \fifo_ram_module/app_addr[12] ;
input \fifo_ram_module/app_addr[11] ;
input \fifo_ram_module/app_addr[10] ;
input \fifo_ram_module/app_addr[9] ;
input \fifo_ram_module/app_addr[8] ;
input \fifo_ram_module/app_addr[7] ;
input \fifo_ram_module/app_addr[6] ;
input \fifo_ram_module/app_addr[5] ;
input \fifo_ram_module/app_addr[4] ;
input \fifo_ram_module/app_addr[3] ;
input \fifo_ram_module/app_addr[2] ;
input \fifo_ram_module/app_addr[1] ;
input \fifo_ram_module/app_addr[0] ;
input \fifo_ram_module/state[3] ;
input \fifo_ram_module/state[2] ;
input \fifo_ram_module/state[1] ;
input \fifo_ram_module/state[0] ;
input \fifo_ram_module/count[31] ;
input \fifo_ram_module/count[30] ;
input \fifo_ram_module/count[29] ;
input \fifo_ram_module/count[28] ;
input \fifo_ram_module/count[27] ;
input \fifo_ram_module/count[26] ;
input \fifo_ram_module/count[25] ;
input \fifo_ram_module/count[24] ;
input \fifo_ram_module/count[23] ;
input \fifo_ram_module/count[22] ;
input \fifo_ram_module/count[21] ;
input \fifo_ram_module/count[20] ;
input \fifo_ram_module/count[19] ;
input \fifo_ram_module/count[18] ;
input \fifo_ram_module/count[17] ;
input \fifo_ram_module/count[16] ;
input \fifo_ram_module/count[15] ;
input \fifo_ram_module/count[14] ;
input \fifo_ram_module/count[13] ;
input \fifo_ram_module/count[12] ;
input \fifo_ram_module/count[11] ;
input \fifo_ram_module/count[10] ;
input \fifo_ram_module/count[9] ;
input \fifo_ram_module/count[8] ;
input \fifo_ram_module/count[7] ;
input \fifo_ram_module/count[6] ;
input \fifo_ram_module/count[5] ;
input \fifo_ram_module/count[4] ;
input \fifo_ram_module/count[3] ;
input \fifo_ram_module/count[2] ;
input \fifo_ram_module/count[1] ;
input \fifo_ram_module/count[0] ;
input \fifo_ram_module/cmd_ready ;
input \fifo_ram_module/cmd_en ;
input \fifo_ram_module/wr_ready ;
input \fifo_ram_module/wr_en ;
input \fifo_ram_module/rd_data_valid ;
input \fifo_ram_module/fifo_read_full ;
input \fifo_ram_module/fifo_write_empty ;
input \fifo_ram_module/fifo_read_almost_empty ;
input \fifo_ram_module/fifo_write_rd_en ;
input \fifo_ram_module/fifo_read_wr_en ;
input \fifo_ram_module/fifo_write_full ;
input \fifo_ram_module/fifo_read_empty ;
input read_en;
input \state[3] ;
input \state[2] ;
input \state[1] ;
input \state[0] ;
input sd_file_found;
input clk;
input tms_pad_i;
input tck_pad_i;
input tdi_pad_i;
output tdo_pad_o;

wire \read_data[15] ;
wire \read_data[14] ;
wire \read_data[13] ;
wire \read_data[12] ;
wire \read_data[11] ;
wire \read_data[10] ;
wire \read_data[9] ;
wire \read_data[8] ;
wire \read_data[7] ;
wire \read_data[6] ;
wire \read_data[5] ;
wire \read_data[4] ;
wire \read_data[3] ;
wire \read_data[2] ;
wire \read_data[1] ;
wire \read_data[0] ;
wire \fifo_ram_module/rd_data[255] ;
wire \fifo_ram_module/rd_data[254] ;
wire \fifo_ram_module/rd_data[253] ;
wire \fifo_ram_module/rd_data[252] ;
wire \fifo_ram_module/rd_data[251] ;
wire \fifo_ram_module/rd_data[250] ;
wire \fifo_ram_module/rd_data[249] ;
wire \fifo_ram_module/rd_data[248] ;
wire \fifo_ram_module/rd_data[247] ;
wire \fifo_ram_module/rd_data[246] ;
wire \fifo_ram_module/rd_data[245] ;
wire \fifo_ram_module/rd_data[244] ;
wire \fifo_ram_module/rd_data[243] ;
wire \fifo_ram_module/rd_data[242] ;
wire \fifo_ram_module/rd_data[241] ;
wire \fifo_ram_module/rd_data[240] ;
wire \fifo_ram_module/rd_data[239] ;
wire \fifo_ram_module/rd_data[238] ;
wire \fifo_ram_module/rd_data[237] ;
wire \fifo_ram_module/rd_data[236] ;
wire \fifo_ram_module/rd_data[235] ;
wire \fifo_ram_module/rd_data[234] ;
wire \fifo_ram_module/rd_data[233] ;
wire \fifo_ram_module/rd_data[232] ;
wire \fifo_ram_module/rd_data[231] ;
wire \fifo_ram_module/rd_data[230] ;
wire \fifo_ram_module/rd_data[229] ;
wire \fifo_ram_module/rd_data[228] ;
wire \fifo_ram_module/rd_data[227] ;
wire \fifo_ram_module/rd_data[226] ;
wire \fifo_ram_module/rd_data[225] ;
wire \fifo_ram_module/rd_data[224] ;
wire \fifo_ram_module/rd_data[223] ;
wire \fifo_ram_module/rd_data[222] ;
wire \fifo_ram_module/rd_data[221] ;
wire \fifo_ram_module/rd_data[220] ;
wire \fifo_ram_module/rd_data[219] ;
wire \fifo_ram_module/rd_data[218] ;
wire \fifo_ram_module/rd_data[217] ;
wire \fifo_ram_module/rd_data[216] ;
wire \fifo_ram_module/rd_data[215] ;
wire \fifo_ram_module/rd_data[214] ;
wire \fifo_ram_module/rd_data[213] ;
wire \fifo_ram_module/rd_data[212] ;
wire \fifo_ram_module/rd_data[211] ;
wire \fifo_ram_module/rd_data[210] ;
wire \fifo_ram_module/rd_data[209] ;
wire \fifo_ram_module/rd_data[208] ;
wire \fifo_ram_module/rd_data[207] ;
wire \fifo_ram_module/rd_data[206] ;
wire \fifo_ram_module/rd_data[205] ;
wire \fifo_ram_module/rd_data[204] ;
wire \fifo_ram_module/rd_data[203] ;
wire \fifo_ram_module/rd_data[202] ;
wire \fifo_ram_module/rd_data[201] ;
wire \fifo_ram_module/rd_data[200] ;
wire \fifo_ram_module/rd_data[199] ;
wire \fifo_ram_module/rd_data[198] ;
wire \fifo_ram_module/rd_data[197] ;
wire \fifo_ram_module/rd_data[196] ;
wire \fifo_ram_module/rd_data[195] ;
wire \fifo_ram_module/rd_data[194] ;
wire \fifo_ram_module/rd_data[193] ;
wire \fifo_ram_module/rd_data[192] ;
wire \fifo_ram_module/rd_data[191] ;
wire \fifo_ram_module/rd_data[190] ;
wire \fifo_ram_module/rd_data[189] ;
wire \fifo_ram_module/rd_data[188] ;
wire \fifo_ram_module/rd_data[187] ;
wire \fifo_ram_module/rd_data[186] ;
wire \fifo_ram_module/rd_data[185] ;
wire \fifo_ram_module/rd_data[184] ;
wire \fifo_ram_module/rd_data[183] ;
wire \fifo_ram_module/rd_data[182] ;
wire \fifo_ram_module/rd_data[181] ;
wire \fifo_ram_module/rd_data[180] ;
wire \fifo_ram_module/rd_data[179] ;
wire \fifo_ram_module/rd_data[178] ;
wire \fifo_ram_module/rd_data[177] ;
wire \fifo_ram_module/rd_data[176] ;
wire \fifo_ram_module/rd_data[175] ;
wire \fifo_ram_module/rd_data[174] ;
wire \fifo_ram_module/rd_data[173] ;
wire \fifo_ram_module/rd_data[172] ;
wire \fifo_ram_module/rd_data[171] ;
wire \fifo_ram_module/rd_data[170] ;
wire \fifo_ram_module/rd_data[169] ;
wire \fifo_ram_module/rd_data[168] ;
wire \fifo_ram_module/rd_data[167] ;
wire \fifo_ram_module/rd_data[166] ;
wire \fifo_ram_module/rd_data[165] ;
wire \fifo_ram_module/rd_data[164] ;
wire \fifo_ram_module/rd_data[163] ;
wire \fifo_ram_module/rd_data[162] ;
wire \fifo_ram_module/rd_data[161] ;
wire \fifo_ram_module/rd_data[160] ;
wire \fifo_ram_module/rd_data[159] ;
wire \fifo_ram_module/rd_data[158] ;
wire \fifo_ram_module/rd_data[157] ;
wire \fifo_ram_module/rd_data[156] ;
wire \fifo_ram_module/rd_data[155] ;
wire \fifo_ram_module/rd_data[154] ;
wire \fifo_ram_module/rd_data[153] ;
wire \fifo_ram_module/rd_data[152] ;
wire \fifo_ram_module/rd_data[151] ;
wire \fifo_ram_module/rd_data[150] ;
wire \fifo_ram_module/rd_data[149] ;
wire \fifo_ram_module/rd_data[148] ;
wire \fifo_ram_module/rd_data[147] ;
wire \fifo_ram_module/rd_data[146] ;
wire \fifo_ram_module/rd_data[145] ;
wire \fifo_ram_module/rd_data[144] ;
wire \fifo_ram_module/rd_data[143] ;
wire \fifo_ram_module/rd_data[142] ;
wire \fifo_ram_module/rd_data[141] ;
wire \fifo_ram_module/rd_data[140] ;
wire \fifo_ram_module/rd_data[139] ;
wire \fifo_ram_module/rd_data[138] ;
wire \fifo_ram_module/rd_data[137] ;
wire \fifo_ram_module/rd_data[136] ;
wire \fifo_ram_module/rd_data[135] ;
wire \fifo_ram_module/rd_data[134] ;
wire \fifo_ram_module/rd_data[133] ;
wire \fifo_ram_module/rd_data[132] ;
wire \fifo_ram_module/rd_data[131] ;
wire \fifo_ram_module/rd_data[130] ;
wire \fifo_ram_module/rd_data[129] ;
wire \fifo_ram_module/rd_data[128] ;
wire \fifo_ram_module/rd_data[127] ;
wire \fifo_ram_module/rd_data[126] ;
wire \fifo_ram_module/rd_data[125] ;
wire \fifo_ram_module/rd_data[124] ;
wire \fifo_ram_module/rd_data[123] ;
wire \fifo_ram_module/rd_data[122] ;
wire \fifo_ram_module/rd_data[121] ;
wire \fifo_ram_module/rd_data[120] ;
wire \fifo_ram_module/rd_data[119] ;
wire \fifo_ram_module/rd_data[118] ;
wire \fifo_ram_module/rd_data[117] ;
wire \fifo_ram_module/rd_data[116] ;
wire \fifo_ram_module/rd_data[115] ;
wire \fifo_ram_module/rd_data[114] ;
wire \fifo_ram_module/rd_data[113] ;
wire \fifo_ram_module/rd_data[112] ;
wire \fifo_ram_module/rd_data[111] ;
wire \fifo_ram_module/rd_data[110] ;
wire \fifo_ram_module/rd_data[109] ;
wire \fifo_ram_module/rd_data[108] ;
wire \fifo_ram_module/rd_data[107] ;
wire \fifo_ram_module/rd_data[106] ;
wire \fifo_ram_module/rd_data[105] ;
wire \fifo_ram_module/rd_data[104] ;
wire \fifo_ram_module/rd_data[103] ;
wire \fifo_ram_module/rd_data[102] ;
wire \fifo_ram_module/rd_data[101] ;
wire \fifo_ram_module/rd_data[100] ;
wire \fifo_ram_module/rd_data[99] ;
wire \fifo_ram_module/rd_data[98] ;
wire \fifo_ram_module/rd_data[97] ;
wire \fifo_ram_module/rd_data[96] ;
wire \fifo_ram_module/rd_data[95] ;
wire \fifo_ram_module/rd_data[94] ;
wire \fifo_ram_module/rd_data[93] ;
wire \fifo_ram_module/rd_data[92] ;
wire \fifo_ram_module/rd_data[91] ;
wire \fifo_ram_module/rd_data[90] ;
wire \fifo_ram_module/rd_data[89] ;
wire \fifo_ram_module/rd_data[88] ;
wire \fifo_ram_module/rd_data[87] ;
wire \fifo_ram_module/rd_data[86] ;
wire \fifo_ram_module/rd_data[85] ;
wire \fifo_ram_module/rd_data[84] ;
wire \fifo_ram_module/rd_data[83] ;
wire \fifo_ram_module/rd_data[82] ;
wire \fifo_ram_module/rd_data[81] ;
wire \fifo_ram_module/rd_data[80] ;
wire \fifo_ram_module/rd_data[79] ;
wire \fifo_ram_module/rd_data[78] ;
wire \fifo_ram_module/rd_data[77] ;
wire \fifo_ram_module/rd_data[76] ;
wire \fifo_ram_module/rd_data[75] ;
wire \fifo_ram_module/rd_data[74] ;
wire \fifo_ram_module/rd_data[73] ;
wire \fifo_ram_module/rd_data[72] ;
wire \fifo_ram_module/rd_data[71] ;
wire \fifo_ram_module/rd_data[70] ;
wire \fifo_ram_module/rd_data[69] ;
wire \fifo_ram_module/rd_data[68] ;
wire \fifo_ram_module/rd_data[67] ;
wire \fifo_ram_module/rd_data[66] ;
wire \fifo_ram_module/rd_data[65] ;
wire \fifo_ram_module/rd_data[64] ;
wire \fifo_ram_module/rd_data[63] ;
wire \fifo_ram_module/rd_data[62] ;
wire \fifo_ram_module/rd_data[61] ;
wire \fifo_ram_module/rd_data[60] ;
wire \fifo_ram_module/rd_data[59] ;
wire \fifo_ram_module/rd_data[58] ;
wire \fifo_ram_module/rd_data[57] ;
wire \fifo_ram_module/rd_data[56] ;
wire \fifo_ram_module/rd_data[55] ;
wire \fifo_ram_module/rd_data[54] ;
wire \fifo_ram_module/rd_data[53] ;
wire \fifo_ram_module/rd_data[52] ;
wire \fifo_ram_module/rd_data[51] ;
wire \fifo_ram_module/rd_data[50] ;
wire \fifo_ram_module/rd_data[49] ;
wire \fifo_ram_module/rd_data[48] ;
wire \fifo_ram_module/rd_data[47] ;
wire \fifo_ram_module/rd_data[46] ;
wire \fifo_ram_module/rd_data[45] ;
wire \fifo_ram_module/rd_data[44] ;
wire \fifo_ram_module/rd_data[43] ;
wire \fifo_ram_module/rd_data[42] ;
wire \fifo_ram_module/rd_data[41] ;
wire \fifo_ram_module/rd_data[40] ;
wire \fifo_ram_module/rd_data[39] ;
wire \fifo_ram_module/rd_data[38] ;
wire \fifo_ram_module/rd_data[37] ;
wire \fifo_ram_module/rd_data[36] ;
wire \fifo_ram_module/rd_data[35] ;
wire \fifo_ram_module/rd_data[34] ;
wire \fifo_ram_module/rd_data[33] ;
wire \fifo_ram_module/rd_data[32] ;
wire \fifo_ram_module/rd_data[31] ;
wire \fifo_ram_module/rd_data[30] ;
wire \fifo_ram_module/rd_data[29] ;
wire \fifo_ram_module/rd_data[28] ;
wire \fifo_ram_module/rd_data[27] ;
wire \fifo_ram_module/rd_data[26] ;
wire \fifo_ram_module/rd_data[25] ;
wire \fifo_ram_module/rd_data[24] ;
wire \fifo_ram_module/rd_data[23] ;
wire \fifo_ram_module/rd_data[22] ;
wire \fifo_ram_module/rd_data[21] ;
wire \fifo_ram_module/rd_data[20] ;
wire \fifo_ram_module/rd_data[19] ;
wire \fifo_ram_module/rd_data[18] ;
wire \fifo_ram_module/rd_data[17] ;
wire \fifo_ram_module/rd_data[16] ;
wire \fifo_ram_module/rd_data[15] ;
wire \fifo_ram_module/rd_data[14] ;
wire \fifo_ram_module/rd_data[13] ;
wire \fifo_ram_module/rd_data[12] ;
wire \fifo_ram_module/rd_data[11] ;
wire \fifo_ram_module/rd_data[10] ;
wire \fifo_ram_module/rd_data[9] ;
wire \fifo_ram_module/rd_data[8] ;
wire \fifo_ram_module/rd_data[7] ;
wire \fifo_ram_module/rd_data[6] ;
wire \fifo_ram_module/rd_data[5] ;
wire \fifo_ram_module/rd_data[4] ;
wire \fifo_ram_module/rd_data[3] ;
wire \fifo_ram_module/rd_data[2] ;
wire \fifo_ram_module/rd_data[1] ;
wire \fifo_ram_module/rd_data[0] ;
wire \fifo_ram_module/cmd[2] ;
wire \fifo_ram_module/cmd[1] ;
wire \fifo_ram_module/cmd[0] ;
wire \fifo_ram_module/app_addr[28] ;
wire \fifo_ram_module/app_addr[27] ;
wire \fifo_ram_module/app_addr[26] ;
wire \fifo_ram_module/app_addr[25] ;
wire \fifo_ram_module/app_addr[24] ;
wire \fifo_ram_module/app_addr[23] ;
wire \fifo_ram_module/app_addr[22] ;
wire \fifo_ram_module/app_addr[21] ;
wire \fifo_ram_module/app_addr[20] ;
wire \fifo_ram_module/app_addr[19] ;
wire \fifo_ram_module/app_addr[18] ;
wire \fifo_ram_module/app_addr[17] ;
wire \fifo_ram_module/app_addr[16] ;
wire \fifo_ram_module/app_addr[15] ;
wire \fifo_ram_module/app_addr[14] ;
wire \fifo_ram_module/app_addr[13] ;
wire \fifo_ram_module/app_addr[12] ;
wire \fifo_ram_module/app_addr[11] ;
wire \fifo_ram_module/app_addr[10] ;
wire \fifo_ram_module/app_addr[9] ;
wire \fifo_ram_module/app_addr[8] ;
wire \fifo_ram_module/app_addr[7] ;
wire \fifo_ram_module/app_addr[6] ;
wire \fifo_ram_module/app_addr[5] ;
wire \fifo_ram_module/app_addr[4] ;
wire \fifo_ram_module/app_addr[3] ;
wire \fifo_ram_module/app_addr[2] ;
wire \fifo_ram_module/app_addr[1] ;
wire \fifo_ram_module/app_addr[0] ;
wire \fifo_ram_module/state[3] ;
wire \fifo_ram_module/state[2] ;
wire \fifo_ram_module/state[1] ;
wire \fifo_ram_module/state[0] ;
wire \fifo_ram_module/count[31] ;
wire \fifo_ram_module/count[30] ;
wire \fifo_ram_module/count[29] ;
wire \fifo_ram_module/count[28] ;
wire \fifo_ram_module/count[27] ;
wire \fifo_ram_module/count[26] ;
wire \fifo_ram_module/count[25] ;
wire \fifo_ram_module/count[24] ;
wire \fifo_ram_module/count[23] ;
wire \fifo_ram_module/count[22] ;
wire \fifo_ram_module/count[21] ;
wire \fifo_ram_module/count[20] ;
wire \fifo_ram_module/count[19] ;
wire \fifo_ram_module/count[18] ;
wire \fifo_ram_module/count[17] ;
wire \fifo_ram_module/count[16] ;
wire \fifo_ram_module/count[15] ;
wire \fifo_ram_module/count[14] ;
wire \fifo_ram_module/count[13] ;
wire \fifo_ram_module/count[12] ;
wire \fifo_ram_module/count[11] ;
wire \fifo_ram_module/count[10] ;
wire \fifo_ram_module/count[9] ;
wire \fifo_ram_module/count[8] ;
wire \fifo_ram_module/count[7] ;
wire \fifo_ram_module/count[6] ;
wire \fifo_ram_module/count[5] ;
wire \fifo_ram_module/count[4] ;
wire \fifo_ram_module/count[3] ;
wire \fifo_ram_module/count[2] ;
wire \fifo_ram_module/count[1] ;
wire \fifo_ram_module/count[0] ;
wire \fifo_ram_module/cmd_ready ;
wire \fifo_ram_module/cmd_en ;
wire \fifo_ram_module/wr_ready ;
wire \fifo_ram_module/wr_en ;
wire \fifo_ram_module/rd_data_valid ;
wire \fifo_ram_module/fifo_read_full ;
wire \fifo_ram_module/fifo_write_empty ;
wire \fifo_ram_module/fifo_read_almost_empty ;
wire \fifo_ram_module/fifo_write_rd_en ;
wire \fifo_ram_module/fifo_read_wr_en ;
wire \fifo_ram_module/fifo_write_full ;
wire \fifo_ram_module/fifo_read_empty ;
wire read_en;
wire \state[3] ;
wire \state[2] ;
wire \state[1] ;
wire \state[0] ;
wire sd_file_found;
wire clk;
wire tms_pad_i;
wire tck_pad_i;
wire tdi_pad_i;
wire tdo_pad_o;
wire tms_i_c;
wire tck_i_c;
wire tdi_i_c;
wire tdo_o_c;
wire [9:0] control0;
wire gao_jtag_tck;
wire gao_jtag_reset;
wire run_test_idle_er1;
wire run_test_idle_er2;
wire shift_dr_capture_dr;
wire update_dr;
wire pause_dr;
wire enable_er1;
wire enable_er2;
wire gao_jtag_tdi;
wire tdo_er1;

IBUF tms_ibuf (
    .I(tms_pad_i),
    .O(tms_i_c)
);

IBUF tck_ibuf (
    .I(tck_pad_i),
    .O(tck_i_c)
);

IBUF tdi_ibuf (
    .I(tdi_pad_i),
    .O(tdi_i_c)
);

OBUF tdo_obuf (
    .I(tdo_o_c),
    .O(tdo_pad_o)
);

GW_JTAG  u_gw_jtag(
    .tms_pad_i(tms_i_c),
    .tck_pad_i(tck_i_c),
    .tdi_pad_i(tdi_i_c),
    .tdo_pad_o(tdo_o_c),
    .tck_o(gao_jtag_tck),
    .test_logic_reset_o(gao_jtag_reset),
    .run_test_idle_er1_o(run_test_idle_er1),
    .run_test_idle_er2_o(run_test_idle_er2),
    .shift_dr_capture_dr_o(shift_dr_capture_dr),
    .update_dr_o(update_dr),
    .pause_dr_o(pause_dr),
    .enable_er1_o(enable_er1),
    .enable_er2_o(enable_er2),
    .tdi_o(gao_jtag_tdi),
    .tdo_er1_i(tdo_er1),
    .tdo_er2_i(1'b0)
);

gw_con_top  u_icon_top(
    .tck_i(gao_jtag_tck),
    .tdi_i(gao_jtag_tdi),
    .tdo_o(tdo_er1),
    .rst_i(gao_jtag_reset),
    .control0(control0[9:0]),
    .enable_i(enable_er1),
    .shift_dr_capture_dr_i(shift_dr_capture_dr),
    .update_dr_i(update_dr)
);

ao_top_0  u_la0_top(
    .control(control0[9:0]),
    .trig0_i({\state[3] ,\state[2] ,\state[1] ,\state[0] }),
    .data_i({\read_data[15] ,\read_data[14] ,\read_data[13] ,\read_data[12] ,\read_data[11] ,\read_data[10] ,\read_data[9] ,\read_data[8] ,\read_data[7] ,\read_data[6] ,\read_data[5] ,\read_data[4] ,\read_data[3] ,\read_data[2] ,\read_data[1] ,\read_data[0] ,\fifo_ram_module/rd_data[255] ,\fifo_ram_module/rd_data[254] ,\fifo_ram_module/rd_data[253] ,\fifo_ram_module/rd_data[252] ,\fifo_ram_module/rd_data[251] ,\fifo_ram_module/rd_data[250] ,\fifo_ram_module/rd_data[249] ,\fifo_ram_module/rd_data[248] ,\fifo_ram_module/rd_data[247] ,\fifo_ram_module/rd_data[246] ,\fifo_ram_module/rd_data[245] ,\fifo_ram_module/rd_data[244] ,\fifo_ram_module/rd_data[243] ,\fifo_ram_module/rd_data[242] ,\fifo_ram_module/rd_data[241] ,\fifo_ram_module/rd_data[240] ,\fifo_ram_module/rd_data[239] ,\fifo_ram_module/rd_data[238] ,\fifo_ram_module/rd_data[237] ,\fifo_ram_module/rd_data[236] ,\fifo_ram_module/rd_data[235] ,\fifo_ram_module/rd_data[234] ,\fifo_ram_module/rd_data[233] ,\fifo_ram_module/rd_data[232] ,\fifo_ram_module/rd_data[231] ,\fifo_ram_module/rd_data[230] ,\fifo_ram_module/rd_data[229] ,\fifo_ram_module/rd_data[228] ,\fifo_ram_module/rd_data[227] ,\fifo_ram_module/rd_data[226] ,\fifo_ram_module/rd_data[225] ,\fifo_ram_module/rd_data[224] ,\fifo_ram_module/rd_data[223] ,\fifo_ram_module/rd_data[222] ,\fifo_ram_module/rd_data[221] ,\fifo_ram_module/rd_data[220] ,\fifo_ram_module/rd_data[219] ,\fifo_ram_module/rd_data[218] ,\fifo_ram_module/rd_data[217] ,\fifo_ram_module/rd_data[216] ,\fifo_ram_module/rd_data[215] ,\fifo_ram_module/rd_data[214] ,\fifo_ram_module/rd_data[213] ,\fifo_ram_module/rd_data[212] ,\fifo_ram_module/rd_data[211] ,\fifo_ram_module/rd_data[210] ,\fifo_ram_module/rd_data[209] ,\fifo_ram_module/rd_data[208] ,\fifo_ram_module/rd_data[207] ,\fifo_ram_module/rd_data[206] ,\fifo_ram_module/rd_data[205] ,\fifo_ram_module/rd_data[204] ,\fifo_ram_module/rd_data[203] ,\fifo_ram_module/rd_data[202] ,\fifo_ram_module/rd_data[201] ,\fifo_ram_module/rd_data[200] ,\fifo_ram_module/rd_data[199] ,\fifo_ram_module/rd_data[198] ,\fifo_ram_module/rd_data[197] ,\fifo_ram_module/rd_data[196] ,\fifo_ram_module/rd_data[195] ,\fifo_ram_module/rd_data[194] ,\fifo_ram_module/rd_data[193] ,\fifo_ram_module/rd_data[192] ,\fifo_ram_module/rd_data[191] ,\fifo_ram_module/rd_data[190] ,\fifo_ram_module/rd_data[189] ,\fifo_ram_module/rd_data[188] ,\fifo_ram_module/rd_data[187] ,\fifo_ram_module/rd_data[186] ,\fifo_ram_module/rd_data[185] ,\fifo_ram_module/rd_data[184] ,\fifo_ram_module/rd_data[183] ,\fifo_ram_module/rd_data[182] ,\fifo_ram_module/rd_data[181] ,\fifo_ram_module/rd_data[180] ,\fifo_ram_module/rd_data[179] ,\fifo_ram_module/rd_data[178] ,\fifo_ram_module/rd_data[177] ,\fifo_ram_module/rd_data[176] ,\fifo_ram_module/rd_data[175] ,\fifo_ram_module/rd_data[174] ,\fifo_ram_module/rd_data[173] ,\fifo_ram_module/rd_data[172] ,\fifo_ram_module/rd_data[171] ,\fifo_ram_module/rd_data[170] ,\fifo_ram_module/rd_data[169] ,\fifo_ram_module/rd_data[168] ,\fifo_ram_module/rd_data[167] ,\fifo_ram_module/rd_data[166] ,\fifo_ram_module/rd_data[165] ,\fifo_ram_module/rd_data[164] ,\fifo_ram_module/rd_data[163] ,\fifo_ram_module/rd_data[162] ,\fifo_ram_module/rd_data[161] ,\fifo_ram_module/rd_data[160] ,\fifo_ram_module/rd_data[159] ,\fifo_ram_module/rd_data[158] ,\fifo_ram_module/rd_data[157] ,\fifo_ram_module/rd_data[156] ,\fifo_ram_module/rd_data[155] ,\fifo_ram_module/rd_data[154] ,\fifo_ram_module/rd_data[153] ,\fifo_ram_module/rd_data[152] ,\fifo_ram_module/rd_data[151] ,\fifo_ram_module/rd_data[150] ,\fifo_ram_module/rd_data[149] ,\fifo_ram_module/rd_data[148] ,\fifo_ram_module/rd_data[147] ,\fifo_ram_module/rd_data[146] ,\fifo_ram_module/rd_data[145] ,\fifo_ram_module/rd_data[144] ,\fifo_ram_module/rd_data[143] ,\fifo_ram_module/rd_data[142] ,\fifo_ram_module/rd_data[141] ,\fifo_ram_module/rd_data[140] ,\fifo_ram_module/rd_data[139] ,\fifo_ram_module/rd_data[138] ,\fifo_ram_module/rd_data[137] ,\fifo_ram_module/rd_data[136] ,\fifo_ram_module/rd_data[135] ,\fifo_ram_module/rd_data[134] ,\fifo_ram_module/rd_data[133] ,\fifo_ram_module/rd_data[132] ,\fifo_ram_module/rd_data[131] ,\fifo_ram_module/rd_data[130] ,\fifo_ram_module/rd_data[129] ,\fifo_ram_module/rd_data[128] ,\fifo_ram_module/rd_data[127] ,\fifo_ram_module/rd_data[126] ,\fifo_ram_module/rd_data[125] ,\fifo_ram_module/rd_data[124] ,\fifo_ram_module/rd_data[123] ,\fifo_ram_module/rd_data[122] ,\fifo_ram_module/rd_data[121] ,\fifo_ram_module/rd_data[120] ,\fifo_ram_module/rd_data[119] ,\fifo_ram_module/rd_data[118] ,\fifo_ram_module/rd_data[117] ,\fifo_ram_module/rd_data[116] ,\fifo_ram_module/rd_data[115] ,\fifo_ram_module/rd_data[114] ,\fifo_ram_module/rd_data[113] ,\fifo_ram_module/rd_data[112] ,\fifo_ram_module/rd_data[111] ,\fifo_ram_module/rd_data[110] ,\fifo_ram_module/rd_data[109] ,\fifo_ram_module/rd_data[108] ,\fifo_ram_module/rd_data[107] ,\fifo_ram_module/rd_data[106] ,\fifo_ram_module/rd_data[105] ,\fifo_ram_module/rd_data[104] ,\fifo_ram_module/rd_data[103] ,\fifo_ram_module/rd_data[102] ,\fifo_ram_module/rd_data[101] ,\fifo_ram_module/rd_data[100] ,\fifo_ram_module/rd_data[99] ,\fifo_ram_module/rd_data[98] ,\fifo_ram_module/rd_data[97] ,\fifo_ram_module/rd_data[96] ,\fifo_ram_module/rd_data[95] ,\fifo_ram_module/rd_data[94] ,\fifo_ram_module/rd_data[93] ,\fifo_ram_module/rd_data[92] ,\fifo_ram_module/rd_data[91] ,\fifo_ram_module/rd_data[90] ,\fifo_ram_module/rd_data[89] ,\fifo_ram_module/rd_data[88] ,\fifo_ram_module/rd_data[87] ,\fifo_ram_module/rd_data[86] ,\fifo_ram_module/rd_data[85] ,\fifo_ram_module/rd_data[84] ,\fifo_ram_module/rd_data[83] ,\fifo_ram_module/rd_data[82] ,\fifo_ram_module/rd_data[81] ,\fifo_ram_module/rd_data[80] ,\fifo_ram_module/rd_data[79] ,\fifo_ram_module/rd_data[78] ,\fifo_ram_module/rd_data[77] ,\fifo_ram_module/rd_data[76] ,\fifo_ram_module/rd_data[75] ,\fifo_ram_module/rd_data[74] ,\fifo_ram_module/rd_data[73] ,\fifo_ram_module/rd_data[72] ,\fifo_ram_module/rd_data[71] ,\fifo_ram_module/rd_data[70] ,\fifo_ram_module/rd_data[69] ,\fifo_ram_module/rd_data[68] ,\fifo_ram_module/rd_data[67] ,\fifo_ram_module/rd_data[66] ,\fifo_ram_module/rd_data[65] ,\fifo_ram_module/rd_data[64] ,\fifo_ram_module/rd_data[63] ,\fifo_ram_module/rd_data[62] ,\fifo_ram_module/rd_data[61] ,\fifo_ram_module/rd_data[60] ,\fifo_ram_module/rd_data[59] ,\fifo_ram_module/rd_data[58] ,\fifo_ram_module/rd_data[57] ,\fifo_ram_module/rd_data[56] ,\fifo_ram_module/rd_data[55] ,\fifo_ram_module/rd_data[54] ,\fifo_ram_module/rd_data[53] ,\fifo_ram_module/rd_data[52] ,\fifo_ram_module/rd_data[51] ,\fifo_ram_module/rd_data[50] ,\fifo_ram_module/rd_data[49] ,\fifo_ram_module/rd_data[48] ,\fifo_ram_module/rd_data[47] ,\fifo_ram_module/rd_data[46] ,\fifo_ram_module/rd_data[45] ,\fifo_ram_module/rd_data[44] ,\fifo_ram_module/rd_data[43] ,\fifo_ram_module/rd_data[42] ,\fifo_ram_module/rd_data[41] ,\fifo_ram_module/rd_data[40] ,\fifo_ram_module/rd_data[39] ,\fifo_ram_module/rd_data[38] ,\fifo_ram_module/rd_data[37] ,\fifo_ram_module/rd_data[36] ,\fifo_ram_module/rd_data[35] ,\fifo_ram_module/rd_data[34] ,\fifo_ram_module/rd_data[33] ,\fifo_ram_module/rd_data[32] ,\fifo_ram_module/rd_data[31] ,\fifo_ram_module/rd_data[30] ,\fifo_ram_module/rd_data[29] ,\fifo_ram_module/rd_data[28] ,\fifo_ram_module/rd_data[27] ,\fifo_ram_module/rd_data[26] ,\fifo_ram_module/rd_data[25] ,\fifo_ram_module/rd_data[24] ,\fifo_ram_module/rd_data[23] ,\fifo_ram_module/rd_data[22] ,\fifo_ram_module/rd_data[21] ,\fifo_ram_module/rd_data[20] ,\fifo_ram_module/rd_data[19] ,\fifo_ram_module/rd_data[18] ,\fifo_ram_module/rd_data[17] ,\fifo_ram_module/rd_data[16] ,\fifo_ram_module/rd_data[15] ,\fifo_ram_module/rd_data[14] ,\fifo_ram_module/rd_data[13] ,\fifo_ram_module/rd_data[12] ,\fifo_ram_module/rd_data[11] ,\fifo_ram_module/rd_data[10] ,\fifo_ram_module/rd_data[9] ,\fifo_ram_module/rd_data[8] ,\fifo_ram_module/rd_data[7] ,\fifo_ram_module/rd_data[6] ,\fifo_ram_module/rd_data[5] ,\fifo_ram_module/rd_data[4] ,\fifo_ram_module/rd_data[3] ,\fifo_ram_module/rd_data[2] ,\fifo_ram_module/rd_data[1] ,\fifo_ram_module/rd_data[0] ,\fifo_ram_module/cmd[2] ,\fifo_ram_module/cmd[1] ,\fifo_ram_module/cmd[0] ,\fifo_ram_module/app_addr[28] ,\fifo_ram_module/app_addr[27] ,\fifo_ram_module/app_addr[26] ,\fifo_ram_module/app_addr[25] ,\fifo_ram_module/app_addr[24] ,\fifo_ram_module/app_addr[23] ,\fifo_ram_module/app_addr[22] ,\fifo_ram_module/app_addr[21] ,\fifo_ram_module/app_addr[20] ,\fifo_ram_module/app_addr[19] ,\fifo_ram_module/app_addr[18] ,\fifo_ram_module/app_addr[17] ,\fifo_ram_module/app_addr[16] ,\fifo_ram_module/app_addr[15] ,\fifo_ram_module/app_addr[14] ,\fifo_ram_module/app_addr[13] ,\fifo_ram_module/app_addr[12] ,\fifo_ram_module/app_addr[11] ,\fifo_ram_module/app_addr[10] ,\fifo_ram_module/app_addr[9] ,\fifo_ram_module/app_addr[8] ,\fifo_ram_module/app_addr[7] ,\fifo_ram_module/app_addr[6] ,\fifo_ram_module/app_addr[5] ,\fifo_ram_module/app_addr[4] ,\fifo_ram_module/app_addr[3] ,\fifo_ram_module/app_addr[2] ,\fifo_ram_module/app_addr[1] ,\fifo_ram_module/app_addr[0] ,\fifo_ram_module/state[3] ,\fifo_ram_module/state[2] ,\fifo_ram_module/state[1] ,\fifo_ram_module/state[0] ,\fifo_ram_module/count[31] ,\fifo_ram_module/count[30] ,\fifo_ram_module/count[29] ,\fifo_ram_module/count[28] ,\fifo_ram_module/count[27] ,\fifo_ram_module/count[26] ,\fifo_ram_module/count[25] ,\fifo_ram_module/count[24] ,\fifo_ram_module/count[23] ,\fifo_ram_module/count[22] ,\fifo_ram_module/count[21] ,\fifo_ram_module/count[20] ,\fifo_ram_module/count[19] ,\fifo_ram_module/count[18] ,\fifo_ram_module/count[17] ,\fifo_ram_module/count[16] ,\fifo_ram_module/count[15] ,\fifo_ram_module/count[14] ,\fifo_ram_module/count[13] ,\fifo_ram_module/count[12] ,\fifo_ram_module/count[11] ,\fifo_ram_module/count[10] ,\fifo_ram_module/count[9] ,\fifo_ram_module/count[8] ,\fifo_ram_module/count[7] ,\fifo_ram_module/count[6] ,\fifo_ram_module/count[5] ,\fifo_ram_module/count[4] ,\fifo_ram_module/count[3] ,\fifo_ram_module/count[2] ,\fifo_ram_module/count[1] ,\fifo_ram_module/count[0] ,\fifo_ram_module/cmd_ready ,\fifo_ram_module/cmd_en ,\fifo_ram_module/wr_ready ,\fifo_ram_module/wr_en ,\fifo_ram_module/rd_data_valid ,\fifo_ram_module/fifo_read_full ,\fifo_ram_module/fifo_write_empty ,\fifo_ram_module/fifo_read_almost_empty ,\fifo_ram_module/fifo_write_rd_en ,\fifo_ram_module/fifo_read_wr_en ,\fifo_ram_module/fifo_write_full ,\fifo_ram_module/fifo_read_empty ,read_en,\state[3] ,\state[2] ,\state[1] ,\state[0] ,sd_file_found}),
    .clk_i(clk)
);

endmodule
